// Description: The purpose of this module is to generate the next shape randomly, using an LFSR

module next_shape(clk, reset, new_block, curr_shape, next_shape);
	input logic		clk, reset, new_block;   //new_block is asserted high when the block
											 //on the playfield reaches the bottom
	
	//curr shape is in playfield, next shape is displayed to the right of playfield
	output logic [2:0] 	curr_shape, next_shape;	
	
	logic [2:0] next_next_shape; 	//random shape generated by LFSR
	logic		q0, q1, q2, d0;

	//LFSR with tag bits 0 and 2 being fed into an XNOR
	//Note: Using XNOR for this application because there are no shape encodings corresponding
	//to 3'b111. XNOR LFSRs cycle through all possibilities except the highest option, where all
	//bits are 1, and are therefore suited to our purpose here
	d_ff dff0(.clk, .reset, .q(q0), .d(d0));
	d_ff dff1(.clk, .reset, .q(q1), .d(q0));
	d_ff dff2(.clk, .reset, .q(q2), .d(q1));
	
	xnor d_in(d0, q0, q2);  //d0 is result of XNOR of q0, q2
	
	assign next_next_shape = {q2, q1, q0};
	
	always_ff @(posedge clk) begin
		if(reset) begin
			curr_shape <= 3'b0;
			next_shape <= 3'b0;
		end
		else if(new_block) begin
			curr_shape <= next_shape;
			next_shape <= next_next_shape;
		end
	end


endmodule 

module next_shape_testbench();
	logic clk, reset, new_block;
	logic [2:0] curr_shape, next_shape;
	
	next_shape dut(.*);
	
	parameter PERIOD = 100;
	
	initial begin
		clk <= 0;
		forever #(PERIOD/2) clk = ~clk;
	end
	
	initial begin
		@(posedge clk);	reset <= 1;
		@(posedge clk);	reset <= 0;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk); new_block <= 1;
		@(posedge clk); new_block <= 0;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);	new_block <= 1;
		@(posedge clk);	new_block <= 0;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		
		$stop();
	
	end
	

endmodule 